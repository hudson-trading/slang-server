module outer;
    module inner;
    endmodule
endmodule
