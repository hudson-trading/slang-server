module test;
    logic foo;
endmodule
