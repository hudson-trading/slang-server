// Intermediate header that includes base definitions
`include "base_defs.svh"

`define MAX_COUNT 256
