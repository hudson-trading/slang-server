`define MY_MACRO value
`define ANOTHER_MACRO
