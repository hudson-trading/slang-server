`define MY_MACRO value

module m;
endmodule
