

`define SOME_MACRO(arg1, arg2) \
  $display("Macro called with %0d and %0d", arg1, arg2); \
  $display("This is a multi-line macro definition.");
