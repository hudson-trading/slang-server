


module Dut  #(
    parameter int a = 0,
    parameter int b = 1
) (
    input logic foo
);


endmodule
