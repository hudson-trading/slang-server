// Base definitions
`define BUS_WIDTH 64
`define ADDR_SIZE 16
