


module tb;
    logic foo;
endmodule
