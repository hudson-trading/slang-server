class MyClass;
    int x;
endclass

class AnotherClass;
endclass
